-- OrCAD Express generated portmap stub file
-- Matches PCB component pinout with simulation model

